`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/10/26 09:51:17
// Design Name: 
// Module Name: ALU_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ALU_test;

    // �ź�����
    reg [31:0] a;
    reg [31:0] b;
    reg [11:0] op;
    wire [31:0] out;

    // ʵ���� ALU ģ��
    ALU myALU(
        .a(a),
        .b(b),
        .op(op),
        .out(out)
    );

    // ��ʼ�������ź�
    initial begin
        a = 32'h00000002; // ������������ a
        b = 32'h00000001; // ������������ b

        // ִ�в�������
        op = 12'b000000000001; // �ӷ�
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b000000000010; // ����
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b000000000100; // �Ƚ� a < b
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b000000001000; // �Ƚ� a < b
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b000000010000; // �߼��� (a | b)
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b000000100000; // �߼��� (a & b)
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b000001000000; // �߼��� (a | b)
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b000010000000; // ��� (a ^ b)
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b000100000000; // �߼����� (a << b[4:0])
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b001000000000; // �߼����� (a >> b[4:0])
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b010000000000; // �������� (a >>> b[4:0])
        #10; // �ȴ� 10 ��ʱ�䵥λ

        op = 12'b100000000000; // �� b ֱ�Ӹ�ֵ�� out
        #10; // �ȴ� 10 ��ʱ�䵥λ

        // ��������Լ�����Ӹ����������

        $finish; // ��������
    end

endmodule

